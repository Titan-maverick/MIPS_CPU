module InstructionMem(
    // 输入信号
    input [31:0] Addr,             // 地址输入，指定从内存中读取的指令的地址

    // 输出信号
    output reg [31:0] Iout         // 指令输出，32位，存储从内存中读取的指令
);

    // 内存存储空间，大小为 129 字节，每个字节为 8 位
    reg [7:0] ram[128:0];          
    integer i;                     // 用于循环初始化内存

    // 读取指令内存时，每次地址变化时执行此块
    always@(Addr)
    begin
        // 初始化一小部分内存（示例数据），根据实际需要，可以加载更多的指令
        ram[0] = 8'b10101000;      // 内存[0]存储 8 位指令数据
        ram[1] = 8'b00000001;      // 内存[1]存储 8 位指令数据
        ram[2] = 8'b00000000;      // 内存[2]存储 8 位指令数据
        ram[3] = 8'b00000000;      // 内存[3]存储 8 位指令数据

        ram[4] = 8'b00100000;      // 内存[4]存储 8 位指令数据
        ram[5] = 8'b00000010;      // 内存[5]存储 8 位指令数据
        ram[6] = 8'b00000000;      // 内存[6]存储 8 位指令数据
        ram[7] = 8'b00000001;      // 内存[7]存储 8 位指令数据

        ram[8] = 8'b00100000;      // 内存[8]存储 8 位指令数据
        ram[9] = 8'b00000011;      // 内存[9]存储 8 位指令数据
        ram[10] = 8'b00000000;     // 内存[10]存储 8 位指令数据
        ram[11] = 8'b00000001;     // 内存[11]存储 8 位指令数据

        ram[12] = 8'b00000000;     // 内存[12]存储 8 位指令数据
        ram[13] = 8'b00100010;     // 内存[13]存储 8 位指令数据
        ram[14] = 8'b00010000;     // 内存[14]存储 8 位指令数据
        ram[15] = 8'b00101101;     // 内存[15]存储 8 位指令数据

        ram[16] = 8'b00000000;     // 内存[16]存储 8 位指令数据
        ram[17] = 8'b00100011;     // 内存[17]存储 8 位指令数据
        ram[18] = 8'b00001000;     // 内存[18]存储 8 位指令数据
        ram[19] = 8'b00100100;     // 内存[19]存储 8 位指令数据

        ram[20] = 8'b00010100;     // 内存[20]存储 8 位指令数据
        ram[21] = 8'b00100011;     // 内存[21]存储 8 位指令数据
        ram[22] = 8'b11111111;     // 内存[22]存储 8 位指令数据
        ram[23] = 8'b11111101;     // 内存[23]存储 8 位指令数据

        ram[24] = 8'b00010000;     // 内存[24]存储 8 位指令数据
        ram[25] = 8'b11000111;     // 内存[25]存储 8 位指令数据
        ram[26] = 8'b11111111;     // 内存[26]存储 8 位指令数据
        ram[27] = 8'b11111001;     // 内存[27]存储 8 位指令数据

        // 读取内存中的 4 个字节，拼接成 32 位指令输出
        Iout[31:24] = ram[Addr];        // 指令的最高 8 位
        Iout[23:16] = ram[Addr+1];      // 指令的次高 8 位
        Iout[15:8] = ram[Addr+2];       // 指令的次低 8 位
        Iout[7:0] = ram[Addr+3];        // 指令的最低 8 位
    end

endmodule
